`timescale 1 ns / 1 ps

//`default_nettype none
`define WIDTH 16

// Modifications for 15kB block ram, and various other modifications
// by IgorM 11-Dec-2017
// Mind the SPI Flash on the UPduino board must be wired as below
// IgorM 13-Jan-2018: removed obsolate HW 
// IgorM 4-Feb-2018: Added 8 interrupts with priority encoder and interrupt's en/dis mask
// IgorM 9-Feb-2018: Added 4x16kWords of Single Port RAM - SPRAM


  // ######   DEFINES for IOs and PERIPHERALs   #################
  
`define addr_pios            16'h8    // 16'h8

`define addr_int_flgs        16'd40   // 
`define addr_int_mask        16'd50   // 

`define addr_ticksl          16'd100  // 
`define addr_ticksh          16'd101  // 
`define addr_tickshh         16'd102  // 

`define addr_tickssl         16'd105  // 
`define addr_tickssh         16'd106  // 
`define addr_ticksshh        16'd107  // 
`define addr_ticksample      16'd109  // 

`define addr_timer1cl        16'd110  // 
`define addr_timer1ch        16'd111  // 

`define addr_porta_in        16'd310  // 
`define addr_porta_out       16'd311  // 
`define addr_porta_dir       16'd312  // 

`define addr_sram_data0       16'd600  // SPRAM 4 x 16kWords large banks
`define addr_sram_data1       16'd601  // 
`define addr_sram_data2       16'd602  // 
`define addr_sram_data3       16'd603  // 
`define addr_sram_addr        16'd610  // 
 
`define addr_uart0           16'h1000 // 16'h1000

`define addr_util1           16'h2000 // 16'h2000


module SB_RAM256x16(
    output wire [15:0] RDATA,
    input  wire RCLK, RCLKE, RE,
    input  wire [7:0] RADDR,
    input  wire WCLK, WCLKE, WE,
    input  wire [7:0] WADDR,
    input  wire [15:0] MASK, WDATA
);
    parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

  wire [15:0] rd;

  SB_RAM40_4K #(
    .WRITE_MODE(0),
    .READ_MODE(0),
    .INIT_0(INIT_0),
    .INIT_1(INIT_1),
    .INIT_2(INIT_2),
    .INIT_3(INIT_3),
    .INIT_4(INIT_4),
    .INIT_5(INIT_5),
    .INIT_6(INIT_6),
    .INIT_7(INIT_7),
    .INIT_8(INIT_8),
    .INIT_9(INIT_9),
    .INIT_A(INIT_A),
    .INIT_B(INIT_B),
    .INIT_C(INIT_C),
    .INIT_D(INIT_D),
    .INIT_E(INIT_E),
    .INIT_F(INIT_F)
  ) _ram1 (
    .RDATA(rd),
    .RADDR(RADDR),
    .RCLK(RCLK), .RCLKE(RCLKE), .RE(RE),
    .WCLK(WCLK), .WCLKE(WCLKE), .WE(WE),
    .WADDR(WADDR),
    .MASK(16'h0000), 
    .WDATA(WDATA) );

  assign RDATA = rd;

endmodule


// @@@@@@@@@@@@@@@@@@@@@@@@@@

module SB_RAM2048x2(
    output wire [1:0] RDATA,
    input  wire RCLK, RCLKE, RE,
    input  wire [10:0] RADDR,
    input  wire WCLK, WCLKE, WE,
    input  wire [10:0] WADDR,
    input  wire [1:0] MASK, WDATA
);
    parameter INIT_0 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_1 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_2 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_3 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_4 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_5 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_6 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_7 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_8 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_9 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
    parameter INIT_F = 256'h0000000000000000000000000000000000000000000000000000000000000000;

  wire [15:0] rd;

  SB_RAM40_4K #(
    .WRITE_MODE(3),
    .READ_MODE(3),
    .INIT_0(INIT_0),
    .INIT_1(INIT_1),
    .INIT_2(INIT_2),
    .INIT_3(INIT_3),
    .INIT_4(INIT_4),
    .INIT_5(INIT_5),
    .INIT_6(INIT_6),
    .INIT_7(INIT_7),
    .INIT_8(INIT_8),
    .INIT_9(INIT_9),
    .INIT_A(INIT_A),
    .INIT_B(INIT_B),
    .INIT_C(INIT_C),
    .INIT_D(INIT_D),
    .INIT_E(INIT_E),
    .INIT_F(INIT_F)
  ) _ram (
    .RDATA(rd),
    .RADDR(RADDR),
    .RCLK(RCLK), .RCLKE(RCLKE), .RE(RE),
    .WCLK(WCLK), .WCLKE(WCLKE), .WE(WE),
    .WADDR(WADDR),
    .MASK(16'h0000), 
    .WDATA({4'b0, WDATA[1], 7'b0, WDATA[0], 3'b0}));

  assign RDATA[0] = rd[3];
  assign RDATA[1] = rd[11];

endmodule

module top(

        input wire oscillator,
        input wire resetq,

        output wire TXD,       // UART TX
        input  wire RXD,       // UART RX

        output wire SPICLK,    // Flash SCK  --- fpga spiclk  pin 15
        input  wire SPISO,     // Flash SDO  --- fpga spisi   pin 17
        output wire SPISI,     // Flash SDI  --- fpga spiso   pin 14
        output wire SPISSB,    // Flash CS   --- fpga spissb  pin 16

        inout wire PORTA0,
        inout wire PORTA1,
        inout wire PORTA2,
        inout wire PORTA3,
        inout wire PORTA4,
        inout wire PORTA5,
        inout wire PORTA6,
        inout wire PORTA7,
        inout wire PORTA8,
        inout wire PORTA9,
        inout wire PORTA10,
        inout wire PORTA11,
        inout wire PORTA12,
        inout wire PORTA13,
        inout wire PORTA14,
        inout wire PORTA15,

        output wire RGB0,
        output wire RGB1,
        output wire RGB2,
 
        input wire INTR0,
        input wire INTR1,
        input wire INTR2,
        input wire INTR3
);

  // ######   CPU CLOCKS   ###################################

   wire clk ;
  
   // ### Option 1: External 30MHz oscillator (3.3V level)
  
   assign clk = oscillator;

   // ### Option 2: Internal PLL based (max 30MHz with IceCube2)
  
   // my_pll my_pll_inst( 
   //                   .REFERENCECLK(oscillator),
   //                   .PLLOUTCORE(clk),
   //                   .PLLOUTGLOBAL(),
   //                   .RESET(1'b1)   );
 
   // ### Option 3: Internal 24MHz (48MHz/2) oscillator
 
   // SB_HFOSC OSCInst0(
   //                  .CLKHFEN(1'b1),
   //                  .CLKHFPU(1'b1),
   //                  .CLKHF(clk)   );
   // defparam OSCInst0.CLKHF_DIV = "0b01";  // 48MHz DIVIDED by 2

  // ######   RAM   ###########################################
  
  wire io_rd, io_wr;
  wire [15:0] mem_addr;
  wire mem_wr;
  wire [15:0] dout;
  wire [15:0] io_din;
  wire [12:0] code_addr;

  reg unlocked = 0;

// Modification for full 15kB of block ram - for the iCE40UP5k
// Includes nucleus.fs from Mecrisp-Ice
// by IgorM, 11 Dec 2017
// fixes IgorM 11 Jan 2018
// fixes IgorM 29 Jan 2018 - (sliteral) fix

wire [15:0] insn0, insn1, insn2, insn3, insn4, insn5, insn6, insn7, insn8;
wire [15:0] insn;

SB_RAM2048x2 #(
                 .INIT_0(256'hb5300f47df9b8224767717b5ef506f6f52f243bdb6324f67f252d3a7427a4b1a),
                 .INIT_1(256'h3b92dd90a698c3c397628142a7c3979a088a67e64199111185670e0c3e7d5b81),
                 .INIT_2(256'hba724ece895f1b1d864c20c5025660ca484b2f0acbe810f0508c465b9c552ab7),
                 .INIT_3(256'h956711c4a0e2dca7c85541e0a797568638c5074a37a24e6f268688888a4281c2),
                 .INIT_4(256'h030a231ad3c382c270f381c341412a4a608a51c90b4a623a79190b0ac3c0054b),
                 .INIT_5(256'h5100520243e2cbab40320338899ac39b4880a2c82b5a7138191801291aca1a80),
                 .INIT_6(256'ha3a9820a2aa048c880db81ea0a3802e302a000280b630a41c0dba8e35383f0e2),
                 .INIT_7(256'h5a6283a3e8aa0213784829434048a2b0bbc23202d0900a0ab8a192ca2b3b4bcb),
                 .INIT_8(256'h301d0a5b426a606a5a5271182903133b5b23082a280383834243480039494039),
                 .INIT_9(256'h89c90448dbf75557694e90995b12c8263a1760431816d09afab221cbf8da5217),
                 .INIT_A(256'hcdbb613d8cc5031fea81cec9b2e8a6c9b8c189ff18035ec11109643d400fc1ed),
                 .INIT_B(256'h109b07878d09aaf2938126662d4fcdc5440d6e0b01d1b985d8ed486b00e909aa),
                 .INIT_C(256'h8c38d545211dc7c3a702ccb51d7c06b988ac8d03b8a485e924b18191acbc020f),
                 .INIT_D(256'h34946543270c596d43ae33033a66212526155bd310120059c24ec4279898a725),
                 .INIT_E(256'h2de697d2f67226a234f70c8dc3d286e6b77f2a3a5e4fdecf09ec1fbf6f7648d2),
                 .INIT_F(256'hcd7152fd05c3991526a17b9d2f5d05a56cddcc940e861d1d2de625804ed68fb6)
             ) _bn00 (
                 .RDATA(insn0[1:0]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[1:0]));

SB_RAM2048x2 #(
                 .INIT_0(256'hcaeb828a8d0928a91b1a1c04aca1819893473aab008590183fca1a13848c9201),
                 .INIT_1(256'h9a5b928ea16937f042a284a801fd02afa52808e8366baca221ebf237116a4898),
                 .INIT_2(256'h4d102311820b88a084e6006617b013a755a3802088209bebc8c80427a4dea0a5),
                 .INIT_3(256'h83bf80c2edcfc0130eb5db4a1b3bd07489c1f67649a0033371349c00eecb1675),
                 .INIT_4(256'h48ca6038a3a30850fafa5168100068e81161805048f01113a8c887198c4cce42),
                 .INIT_5(256'h085a42990000e1f932e24919f89a7302d3c1606079792060302801b3685ae35b),
                 .INIT_6(256'h022002011171420280911010e22b202021a922a248c8200aa8a9116889811830),
                 .INIT_7(256'h2011c1e01961618168300839100070717070da710a1121a111295848c8290141),
                 .INIT_8(256'hc8088a8a026280c19a918ac28b83f098c1d3b89982bb500081118a0a310000d1),
                 .INIT_9(256'hd45444e49c9001809c187c1c0060e8ac29210286840896e550338004111d29c7),
                 .INIT_A(256'h245f0621724b61717e4f635f233747474846526b769e083a6a36262f82670d39),
                 .INIT_B(256'hf40ae4240664011951197723ecbe4526481803464054681c000591458953c667),
                 .INIT_C(256'h1dc93f9da33d3622899d3428031d2515404b571e491b0b357223403c6435a204),
                 .INIT_D(256'h20bad460a1811b99c24b0e9e451583811394a44411f08058a32421d50c05c0cc),
                 .INIT_E(256'h969e09180d5dcb8d84b52ce99b12050106060f40da1a6c743a084c0e20908119),
                 .INIT_F(256'h131b909040488399868048984545c0e492707818919d491de8ee94a4c34b1918)
             ) _bn01 (
                 .RDATA(insn0[3:2]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[3:2]));

SB_RAM2048x2 #(
                 .INIT_0(256'h20048a20004009a5111013e308988a10d020836c01410920d181127400300fa0),
                 .INIT_1(256'hc8942e776010dd0428480560c61e89280d04e90184108b0bc2a84705f90ccf3d),
                 .INIT_2(256'h908804b0e5761a26c22e04c887bc809a47063024690d08d22aba879a55202390),
                 .INIT_3(256'he4260a62f314c9209a9ec1f602105420a95f74a0fd1d36b57140af87c9382e48),
                 .INIT_4(256'h0820b001380830617082014220a2b058a10be02a00208298302aabb1cca40803),
                 .INIT_5(256'h01a1c008806098721221d189120a206942ea30582379608a79c19a0a8248ab29),
                 .INIT_6(256'h3258023870c802f2110a017b4a620071da7a8038094b0b98080271120ab27311),
                 .INIT_7(256'ha00079180800205968c1294a6039330371011040634300413a431079630841a0),
                 .INIT_8(256'h80c700716901c100f05299088042e870ab08e912d25039592a2b988b99c83903),
                 .INIT_9(256'h89699873843059028600211800288ceba4a900039597132a225cb47f8c960a39),
                 .INIT_A(256'h399c5542718a054c60885884246c3479a3495b08a3e101a045076c40a8120896),
                 .INIT_B(256'h23900890072612529888776362204575465b21205898346305204071669322c1),
                 .INIT_C(256'h1e0438a0a0001c3cacb41c491d64278e0a2e23006044a2c0388a3c282c084a03),
                 .INIT_D(256'h0200435dd110939aa85c0a268004a08ca4bbf010584968abd7012d1264c82101),
                 .INIT_E(256'h0446b06cdc840b14394ac854a2960074034acf5012430845216c12b090b1f421),
                 .INIT_F(256'h8ab4002c80ad90440818b32f285465634010ca790a04938e885c131180588bfa)
             ) _bn02 (
                 .RDATA(insn0[5:4]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[5:4]));

SB_RAM2048x2 #(
                 .INIT_0(256'hca00108bc140808b8211080388081090038040c2000190098281486204008b8b),
                 .INIT_1(256'h369c757da1202a260a68ad105f1c2a01a00d02890684448f09ca7043084140c3),
                 .INIT_2(256'h6c0511122220200224260044608403803406842481213b587032a0a780050a23),
                 .INIT_3(256'h634098ca1cd350c19aa00b820902301002d0a25440d7a116a831b0a31611186a),
                 .INIT_4(256'h20286031ab3808f00070200810a13838500020a07008410098087030848883cb),
                 .INIT_5(256'h0081524a114301d2001040d0e81a0380283932302028006040e1610a082a108a),
                 .INIT_6(256'h1012000109d81040801310810040000053da42800003b0abb00a11c1011a0843),
                 .INIT_7(256'h102099701100600060a010004020403900f162104801310000180080084a0013),
                 .INIT_8(256'hef809a000221088158903298498050a840a910a940d269393b28328000914031),
                 .INIT_9(256'hb42834b810945030bf00b4402c204104098420002095a423dc1810b731941120),
                 .INIT_A(256'h9c2060148a517801c640e63013441a3490231042f4a32c211847522c01a9b514),
                 .INIT_B(256'hd463ac08676c130041182170fc8279e4501222011c486817112440109876c522),
                 .INIT_C(256'h455ca77a77a72e28fd576078063332014002554729001b224f7b003c536f3218),
                 .INIT_D(256'h380098c9b091288f6ac027229100e9c00bab04b0095988e02055301dc886e800),
                 .INIT_E(256'h90840c850180c4c9048944ec82a20d0c868a47c71ad3002018090e1221b161f0),
                 .INIT_F(256'h0d0e90800f0f0302888809aa0d2cc2a0028269e89d8e0c8e2c0c828363c80888)
             ) _bn03 (
                 .RDATA(insn0[7:6]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[7:6]));

SB_RAM2048x2 #(
                 .INIT_0(256'h17300020baf8f020355460204e62707c0a22a869bc53e06500a3024148088b23),
                 .INIT_1(256'h8302b0dcadaa00e05419101019940e828c830579060d18943ea14ac00d224060),
                 .INIT_2(256'ha2f59c6ad4a35044b0a2c29a185b11d14080406598aedd9289d800c24226c5d5),
                 .INIT_3(256'h2f4040a001154c481de7d01749c19096482a0406487d095b64b650f680a165a8),
                 .INIT_4(256'h9808ab2800e84213a3e2594a48b26278234a88ea8b4801aa113390b814e450a3),
                 .INIT_5(256'h01a16a482962e13b2831c86822994138d088e8f8d878008a23e82022604280aa),
                 .INIT_6(256'h89fa4179412a0a222888202960383b3b2a78203060c3a00a19d8592888a142a0),
                 .INIT_7(256'hcae0ab3b8080212960a12003d25122b009111a3bb161105909eb4869522b1872),
                 .INIT_8(256'h88be488a10d09ac9d19198b88283c081a88ae1caabc8293b023b10134280c183),
                 .INIT_9(256'h4248687335f05612604a8a883b3b2a225c9dfecb505028ab91ba001c301c8406),
                 .INIT_A(256'h9083440381b2091ee9fac0ab000a49dfe8ec8aa702822062c9095510a68ab8d3),
                 .INIT_B(256'h80e6869764371086280c603084e72272fc1a032a320b0023045041199b9fa882),
                 .INIT_C(256'h62240026a4ba74eb98bc9de9441a407b9801643320a2080b30ca1c1c346a0c16),
                 .INIT_D(256'h55c4980802120249fb1241648c2e2875181e966220bc2d03d0c01c71e0e52326),
                 .INIT_E(256'h43c24115035221f9023e471959fd4ed220c46432143c8080090d8493b7c6d031),
                 .INIT_F(256'h181c56f52b0f217245dd091dca6b52a6345b79194ccb0c1a6f7a4f8d15561c5c)
             ) _bn04 (
                 .RDATA(insn0[9:8]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[9:8]));

SB_RAM2048x2 #(
                 .INIT_0(256'h00920402222222d01013214003a3226080882892001922c10023000102000093),
                 .INIT_1(256'h03ab08a000032a00066412ba020000330b0a1e04049600c82050408282414390),
                 .INIT_2(256'h22eaa28000c000651082124212608005006080720210a061a041002400f58259),
                 .INIT_3(256'h024a0a5001404113062002c2045d02a012e000e444a000b416c4224100a12060),
                 .INIT_4(256'h083a82003b120242b33160b0a08840002311080000308019002100c015073a48),
                 .INIT_5(256'h8183421120082151a008e812321112628020480070800018a0a221426000003a),
                 .INIT_6(256'h080000400243021008102011305320082200a0c0e001a11918090040881000c0),
                 .INIT_7(256'ha07108000030234080c020108200223021631b71304000020312481212400001),
                 .INIT_8(256'h8060c858a002229133fb00a102c800d2008020ba0280384242500020c2502070),
                 .INIT_9(256'h602a400426068ecc808428b20316224180424250b0f4080100c400056060a0b0),
                 .INIT_A(256'h00a6227220f4004500b800d50010452064b802d62262000e06d310400a9d088c),
                 .INIT_B(256'h23a40b8916470420042820700af802500be20123016502eb1808055023e602c0),
                 .INIT_C(256'h127e28b80090083800a011b98080016000111241000a02123236009800080114),
                 .INIT_D(256'h04ec809004252223a0e000c184901808100094900490a1b5089c0c2c44d10009),
                 .INIT_E(256'h6220000b212000080b05084a50414808101000400008000000148818808180c0),
                 .INIT_F(256'h1141055102230020014000054020227230203061014200006020024b11241000)
             ) _bn05 (
                 .RDATA(insn0[11:10]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[11:10]));

SB_RAM2048x2 #(
                 .INIT_0(256'h7f013602330174406f10e10053006c04ab08bf00fb88f5852b008702fe02b000),
                 .INIT_1(256'h2b0428005b0bc00857114216810193012f067d01ab80b088b703aa02a3803100),
                 .INIT_2(256'hb220e9005700c5009a009a801404cf05ca86eb813c10a701a9005e045707d500),
                 .INIT_3(256'h0b0022080f02270065006e00cd000600040007011e005f05560051151300b303),
                 .INIT_4(256'hdb118880d3089300bb01f200fa08c2000b01cb818a00ab808300080473017800),
                 .INIT_5(256'hab00a1002808f980b988ba80b1019a009000c800d800bb21aa00b3006200ca00),
                 .INIT_6(256'he90178406300a800a800eb016b117a0a2900ba00e100ab80e910ba00a108e200),
                 .INIT_7(256'heb89a208a1003b00c100c3008b00f200bb083128b0107b00e302eb003110f901),
                 .INIT_8(256'h9184d900f222730161110200030053022b212b0b2b09b28a51001300ca00e380),
                 .INIT_9(256'h7f024b08ef08c60ceaa43e0013003200df04ffa0e2c48d0123014c00efa0a784),
                 .INIT_A(256'h2320350037053305150148000900e520e400b3042600c303a58137353e206b24),
                 .INIT_B(256'h2b0f37085404e500a5003020df121300a9001b00a300a200de843d0023062e20),
                 .INIT_C(256'h790c3d101810d3088300b102da80f940f50156008700c100b200b526bfa43d2c),
                 .INIT_D(256'hd710908087004121e700c400af8295081600f710b500f7c47c006708d5015600),
                 .INIT_E(256'h73015200730039015f005b005c00f3087400f5000c0083024501bf00d690d100),
                 .INIT_F(256'h71007f002000750055001400730035107d007800530012007b034c4017007e00)
             ) _bn06 (
                 .RDATA(insn0[13:12]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[13:12]));

SB_RAM2048x2 #(
                 .INIT_0(256'h807b50b604f300fc906f04b98057006c44bb00ef00ff1075441b00ff00f64429),
                 .INIT_1(256'h40bb00d800df20c000b2a8c000e960bf50b9007900eb40f000f754aa007b4429),
                 .INIT_2(256'h085600dd081320dd413f00bb207c00ef20ba006a403400bf04d100de802f08dd),
                 .INIT_3(256'h807b15b2807ed02700dd00be00ef69b61084886640b6807d08b220d9402b00bb),
                 .INIT_4(256'h00fa006820d3009300fa00f200ca01ca304a00fa30d2007b00db407800f200b8),
                 .INIT_5(256'h00fb50f1106800bb00f9407a00d9009a00ea01ea20d200ba00fa409b015a10da),
                 .INIT_6(256'h00eb807800bb11e840b810eb803b806a002141ba10e1500900fb00aa40a100b2),
                 .INIT_7(256'h106300f212e1c05b0299b05b00db00f000b3c03000c0806b00e100fb806900e9),
                 .INIT_8(256'h405a20cb08f200f1188000d278d3008300fb10fb00e840928051600b20ca00b3),
                 .INIT_9(256'h905f044b20ff00931069004e8452707a00d700ff104a00df64fa004e00df0047),
                 .INIT_A(256'h04fb883500dfc03b08e604aaa05b00ff186500ebc01d0cdb30fd802600ee00eb),
                 .INIT_B(256'h00cb40b7841000fd0aada034001f04ea20ad906b04ff488202fc822d00e950af),
                 .INIT_C(256'h009980dd409a20c740260ad5807c00df00ed803a08ff10dd04fe4ab500fcc02f),
                 .INIT_D(256'h28df442068a70479009f02d4503f02f5401408e702bc005f006600c7003518e6),
                 .INIT_E(256'h04faa85e807700ffa05f803f22dc00f702f400b8224d44bbb25d40bd08760699),
                 .INIT_F(256'h807d00fed004887d22d8c01c00ff08fd807c861000dfc01e807600f8a8778076)
             ) _bn07 (
                 .RDATA(insn0[15:14]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[15:14]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000101010101010000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn10 (
                 .RDATA(insn1[1:0]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]  & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[1:0]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000101000001000100),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn11 (
                 .RDATA(insn1[3:2]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]  & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[3:2]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000001000001010000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn12 (
                 .RDATA(insn1[5:4]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]  & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[5:4]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000100000001010101),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn13 (
                 .RDATA(insn1[7:6]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]  & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[7:6]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000101000000010001),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn14 (
                 .RDATA(insn1[9:8]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]  & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[9:8]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000001000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn15 (
                 .RDATA(insn1[11:10]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]  & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[11:10]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn16 (
                 .RDATA(insn1[13:12]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]  & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[13:12]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000010000010001),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn17 (
                 .RDATA(insn1[15:14]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & mem_addr[12]  & !mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[15:14]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn20 (
                 .RDATA(insn2[1:0]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[1:0]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn21 (
                 .RDATA(insn2[3:2]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[3:2]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn22 (
                 .RDATA(insn2[5:4]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[5:4]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn23 (
                 .RDATA(insn2[7:6]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[7:6]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn24 (
                 .RDATA(insn2[9:8]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[9:8]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn25 (
                 .RDATA(insn2[11:10]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[11:10]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn26 (
                 .RDATA(insn2[13:12]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[13:12]));

SB_RAM2048x2 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn27 (
                 .RDATA(insn2[15:14]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked), .WE(mem_wr & !mem_addr[12] & mem_addr[13]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000), .WDATA(dout[15:14]));

// ################################


SB_RAM256x16 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn30 (
                 .RDATA(insn3[15:0]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked),
                 .WE(mem_wr & mem_addr[13] & mem_addr[12] & !mem_addr[11] & !mem_addr[10] & !mem_addr[9]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000),
                 .WDATA(dout[15:0]));


SB_RAM256x16 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn31 (
                 .RDATA(insn4[15:0]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked),
                 .WE(mem_wr & mem_addr[13] & mem_addr[12] & !mem_addr[11] & !mem_addr[10] & mem_addr[9]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000),
                 .WDATA(dout[15:0]));


SB_RAM256x16 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn32 (
                 .RDATA(insn5[15:0]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked),
                 .WE(mem_wr & mem_addr[13] & mem_addr[12] & !mem_addr[11] & mem_addr[10] & !mem_addr[9]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000),
                 .WDATA(dout[15:0]));

SB_RAM256x16 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn33 (
                 .RDATA(insn6[15:0]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked),
                 .WE(mem_wr & mem_addr[13] & mem_addr[12] & !mem_addr[11] & mem_addr[10] & mem_addr[9]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000),
                 .WDATA(dout[15:0]));

SB_RAM256x16 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn34 (
                 .RDATA(insn7[15:0]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked),
                 .WE(mem_wr & mem_addr[13] & mem_addr[12] & mem_addr[11] & !mem_addr[10] & !mem_addr[9]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000),
                 .WDATA(dout[15:0]));


SB_RAM256x16 #(
                 .INIT_0(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_1(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_2(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_3(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_4(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_5(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_6(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_7(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_8(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_9(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_A(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_B(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_C(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_D(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_E(256'h0000000000000000000000000000000000000000000000000000000000000000),
                 .INIT_F(256'h0000000000000000000000000000000000000000000000000000000000000000)
             ) _bn35 (
                 .RDATA(insn8[15:0]),
                 .RADDR(code_addr[10:0]),
                 .RCLK(clk), .RCLKE(1'b1), .RE(1'b1),
                 .WCLK(clk), .WCLKE(unlocked),
                 .WE(mem_wr & mem_addr[13] & mem_addr[12] & mem_addr[11] & !mem_addr[10] & mem_addr[9]),
                 .WADDR(mem_addr[11:1]),
                 .MASK(16'h0000),
                 .WDATA(dout[15:0]));


// ##############################

reg c12, c11, c10, c9, c8;
always @(posedge clk)
begin
    {c12, c11, c10, c9, c8} <= {code_addr[12], code_addr[11], code_addr[10], code_addr[9], code_addr[8]};
end

always @*
begin
    insn = 16'bx;
    casez ({c12, c11}) // Depending on memory address, select different RAM blocks.
        2'b00: insn = insn0;
        2'b01: insn = insn1;
        2'b10: insn = insn2;
        2'b11: begin
            if (!c10 & !c9 & !c8) insn = insn3;   // Select the 256x16 blocks
            if (!c10 & !c9 &  c8) insn = insn4;
            if (!c10 &  c9 & !c8) insn = insn5;
            if (!c10 &  c9 &  c8) insn = insn6;
            if ( c10 & !c9 & !c8) insn = insn7;
            if ( c10 & !c9 &  c8) insn = insn8;
        end

    endcase
end




  // ######   j1a CPU   ########################################
  
    reg [7:0] interrupt = 0;       // up to 8 Interrupts pending, the bit 7 is the highest priority interrupt
    reg [7:0] int_mask  = 0;       // intr enable mask - 1 means the x-th interrupt is enabled
    reg [7:0] int_flags = 8'hFF;   // flags for clearing the processed interrupts (off the ISRs)

  j1 _j1(
    .clk(clk),
    .resetq(resetq),
    .io_rd(io_rd),
    .io_wr(io_wr),
    .mem_wr(mem_wr),
    .dout(dout),
    .io_din(io_din),
    .mem_addr(mem_addr),
    .code_addr(code_addr),
    .insn_from_memory(insn),
    .int_rqst( (interrupt & int_mask) )
  );
  

  // ######   INT_0  RISING EDGE  ################################
  
  reg [2:0] int0dly;
  wire int0re;
  
  // INT0 input synchronizer and edge detector
  
    always @(posedge clk) 
        int0dly <= {int0dly[1:0], INTR0};
 
    assign int0re = (int0dly[2:1] == 2'b01);     // rising edge detector
    // assign int0fe = (int0dly[2:1] == 2'b10);  // falling edge detector

    always @(posedge clk)
    if (int0re == 1)
        interrupt[0] <= 1;
    else
        interrupt[0] <= interrupt[0] & int_flags[0];
        
  // ######   INT_1  RISING EDGE  ################################
  
  reg [2:0] int1dly;
  wire int1re;
  
  // INT1 input synchronizer and edge detector
  
    always @(posedge clk) 
        int1dly <= {int1dly[1:0], INTR1};
 
    assign int1re = (int1dly[2:1] == 2'b01);     // rising edge detector
    // assign int1fe = (int1dly[2:1] == 2'b10);  // falling edge detector
    
    always @(posedge clk)
    if (int1re == 1)
        interrupt[1] <= 1;
    else
        interrupt[1] <= interrupt[1] & int_flags[1];

  // ######   INT_2  RISING EDGE  ################################
  
  reg [2:0] int2dly;
  wire int2re;
  
  // INT2 input synchronizer and edge detector
  
    always @(posedge clk) 
        int2dly <= {int2dly[1:0], INTR2};
 
    assign int2re = (int2dly[2:1] == 2'b01);     // rising edge detector
    // assign int2fe = (int2dly[2:1] == 2'b10);  // falling edge detector
 
    always @(posedge clk)
    if (int2re == 1)
        interrupt[2] <= 1;
    else
        interrupt[2] <= interrupt[2] & int_flags[2];

  // ######   INT_3  RISING SEDGE  ################################
  
  reg [2:0] int3dly;
  wire int3re;
  
  // INT3 input synchronizer and edge detector
  
    always @(posedge clk) 
        int3dly <= {int3dly[1:0], INTR3};
 
    assign int3re = (int3dly[2:1] == 2'b01);     // rising edge detector
    // assign int3fe = (int3dly[2:1] == 2'b10);  // falling edge detector
 
    always @(posedge clk)
    if (int3re == 1)
        interrupt[3] <= 1;
    else
        interrupt[3] <= interrupt[3] & int_flags[3];


  // ######   48 bit CPU TICKS   ##################################

  reg  [47:0] ticks = 0;
  reg  [47:0] tickss = 0;

  // timer ticks

  wire [47:0] ticks_plus_1 = ticks + 1;

  always @(posedge clk)
     ticks <= ticks_plus_1;

  // sample the ticks with "now"

  always @(posedge clk)
     if (io_wr & (mem_addr == `addr_ticksample))  tickss[47:0] <= ticks;


  // ###########  Periodic Timer1 (millis) INTERRUPT 7  ########

  reg [31:0] timer1 = 0;
  reg [31:0] timer1c = 0;

  wire [31:0] timer1_minus_1 = timer1 - 1;

  always @(posedge clk)
    if ( (io_wr & (mem_addr == `addr_timer1ch)) || ( interrupt[7] == 1 ) )
        timer1[31:0] <= timer1c[31:0];
    else
        timer1 <= timer1_minus_1;

  always @(posedge clk)                               // Generate interrupt INT_7 on timer1 compare
    if (timer1 == 1) 
        interrupt[7] <= 1;                            // Set the interrupt INT_7
    else
                                                      // Example of clearing the interrupt pending flag:
        interrupt[7] <= interrupt[7] & int_flags[7];  // Clear the pending interrupt (off the ISR)
        

  // ######   PORTA   ###########################################

  reg  [15:0] porta_dir;   // 1:output, 0:input
  reg  [15:0] porta_out;
  wire [15:0] porta_in;

  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa0  (.PACKAGE_PIN(PORTA0),  .D_OUT_0(porta_out[0]),  .D_IN_0(porta_in[0]),  .OUTPUT_ENABLE(porta_dir[0]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa1  (.PACKAGE_PIN(PORTA1),  .D_OUT_0(porta_out[1]),  .D_IN_0(porta_in[1]),  .OUTPUT_ENABLE(porta_dir[1]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa2  (.PACKAGE_PIN(PORTA2),  .D_OUT_0(porta_out[2]),  .D_IN_0(porta_in[2]),  .OUTPUT_ENABLE(porta_dir[2]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa3  (.PACKAGE_PIN(PORTA3),  .D_OUT_0(porta_out[3]),  .D_IN_0(porta_in[3]),  .OUTPUT_ENABLE(porta_dir[3]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa4  (.PACKAGE_PIN(PORTA4),  .D_OUT_0(porta_out[4]),  .D_IN_0(porta_in[4]),  .OUTPUT_ENABLE(porta_dir[4]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa5  (.PACKAGE_PIN(PORTA5),  .D_OUT_0(porta_out[5]),  .D_IN_0(porta_in[5]),  .OUTPUT_ENABLE(porta_dir[5]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa6  (.PACKAGE_PIN(PORTA6),  .D_OUT_0(porta_out[6]),  .D_IN_0(porta_in[6]),  .OUTPUT_ENABLE(porta_dir[6]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa7  (.PACKAGE_PIN(PORTA7),  .D_OUT_0(porta_out[7]),  .D_IN_0(porta_in[7]),  .OUTPUT_ENABLE(porta_dir[7]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa8  (.PACKAGE_PIN(PORTA8),  .D_OUT_0(porta_out[8]),  .D_IN_0(porta_in[8]),  .OUTPUT_ENABLE(porta_dir[8]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa9  (.PACKAGE_PIN(PORTA9),  .D_OUT_0(porta_out[9]),  .D_IN_0(porta_in[9]),  .OUTPUT_ENABLE(porta_dir[9]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa10 (.PACKAGE_PIN(PORTA10), .D_OUT_0(porta_out[10]), .D_IN_0(porta_in[10]), .OUTPUT_ENABLE(porta_dir[10]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa11 (.PACKAGE_PIN(PORTA11), .D_OUT_0(porta_out[11]), .D_IN_0(porta_in[11]), .OUTPUT_ENABLE(porta_dir[11]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa12 (.PACKAGE_PIN(PORTA12), .D_OUT_0(porta_out[12]), .D_IN_0(porta_in[12]), .OUTPUT_ENABLE(porta_dir[12]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa13 (.PACKAGE_PIN(PORTA13), .D_OUT_0(porta_out[13]), .D_IN_0(porta_in[13]), .OUTPUT_ENABLE(porta_dir[13]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa14 (.PACKAGE_PIN(PORTA14), .D_OUT_0(porta_out[14]), .D_IN_0(porta_in[14]), .OUTPUT_ENABLE(porta_dir[14]));
  SB_IO #(.PIN_TYPE(6'b1010_01)) ioa15 (.PACKAGE_PIN(PORTA15), .D_OUT_0(porta_out[15]), .D_IN_0(porta_in[15]), .OUTPUT_ENABLE(porta_dir[15]));  
  

// ######   UART   ##########################################

  // an RxD 3FF input synchroniser

  reg [2:0] rxddly;
  always @(posedge clk)
    rxddly <= {rxddly[1:0], RXD}; 

  wire uart0_valid, uart0_busy;
  wire [7:0] uart0_data;
  wire uart0_wr = io_wr & (mem_addr == `addr_uart0);
  wire uart0_rd = io_rd & (mem_addr == `addr_uart0);
  wire UART0_RX;
  buart _uart0 (
     .clk(clk),
     .resetq(1'b1),
     .rx(rxddly[2]),
     .tx(TXD),
     .rd(uart0_rd),
     .wr(uart0_wr),
     .valid(uart0_valid),
     .busy(uart0_busy),
     .tx_data(dout[7:0]),
     .rx_data(uart0_data));

  // ######  PIOS   ###################################

  reg [2:0] PIOS;
  assign {SPICLK, SPISI, SPISSB} = PIOS;
 
  wire random = 1; 
  

  // ######   IO PORTS   ######################################

 // READ THE IO REGISTERS
 
  assign io_din =
  
    ((mem_addr == `addr_int_flgs)    ?   int_flags           : 16'd0) |
    ((mem_addr == `addr_int_mask)    ?   int_mask            : 16'd0) |
    
    ((mem_addr == `addr_porta_in)    ?   porta_in            : 16'd0) |
    ((mem_addr == `addr_porta_out)   ?   porta_out           : 16'd0) |
    ((mem_addr == `addr_porta_dir)   ?   porta_dir           : 16'd0) |

    ((mem_addr == `addr_pios)        ?   { 13'd0, PIOS}      : 16'd0) |
    
    ((mem_addr == `addr_sram_data0)   ?   sram_in0[15:0]      : 16'd0) |
    ((mem_addr == `addr_sram_data1)   ?   sram_in1[15:0]      : 16'd0) |
    ((mem_addr == `addr_sram_data2)   ?   sram_in2[15:0]      : 16'd0) |
    ((mem_addr == `addr_sram_data3)   ?   sram_in3[15:0]      : 16'd0) |

    ((mem_addr == `addr_uart0)       ?   { 8'd0, uart0_data} : 16'd0) |
    ((mem_addr == `addr_util1)       ?   {10'd0, random, 2'b00, SPISO, uart0_valid, !uart0_busy} : 16'd0) |

    ((mem_addr == `addr_tickssl)     ?   tickss[15:0]        : 16'd0)|
    ((mem_addr == `addr_tickssh)     ?   tickss[31:16]       : 16'd0)|
    ((mem_addr == `addr_ticksshh)    ?   tickss[47:32]       : 16'd0) ;


 // WRITE THE IO REGISTERS
 
  always @(posedge clk) begin
  
    if (io_wr & (mem_addr == `addr_int_flgs))    int_flags <= dout;
    if (io_wr & (mem_addr == `addr_int_mask))    int_mask <= dout;

    if (io_wr & (mem_addr == `addr_porta_out))   porta_out <= dout;
    if (io_wr & (mem_addr == `addr_porta_dir))   porta_dir <= dout;
    
    if (io_wr & (mem_addr == `addr_pios))        {PIOS} <= dout[2:0];

    if (io_wr & (mem_addr == `addr_timer1cl))    timer1c[15:0] <= dout;
    if (io_wr & (mem_addr == `addr_timer1ch))    timer1c[31:16] <= dout;
    
    if (io_wr & (mem_addr == `addr_sram_addr))   sram_addr[15:0] <= dout;

  end

 
  // ######   MEMLOCK   ########################################

  // This is a workaround to protect memory contents during Reset.
  // Somehow it happens sometimes that the first memory location is corrupted during startup,
  // and as an IO write is one of the earliest things which are done, memory write access is unlocked
  // only after the processor is up and running and sending its welcome message.

  always @(negedge resetq or posedge clk)
  if (!resetq) unlocked <= 0;
  else         unlocked <= unlocked | io_wr;
  
  
  // ######   RGB Tx/Rx indicator   ############################

  defparam RGBA_DRIVER.CURRENT_MODE = "0b1";

  defparam RGBA_DRIVER.RGB0_CURRENT = "0b000001";
  defparam RGBA_DRIVER.RGB1_CURRENT = "0b000001";
  defparam RGBA_DRIVER.RGB2_CURRENT = "0b000001";

    SB_RGBA_DRV RGBA_DRIVER (
        .CURREN(1'b1),
        .RGBLEDEN(1'b1),
        .RGB0PWM(~TXD),
        .RGB1PWM(~RXD),
        .RGB2PWM(0),
        .RGB0(RGB0),
        .RGB1(RGB1),
        .RGB2(RGB2)
    );
    

  // ######  4 x 16kW SPRAM  - Single Port RAM   #################
  
  reg  [15:0] sram_addr;
  
  wire [15:0] sram_in0;
  reg  [15:0] sram_out0;
  
  wire [15:0] sram_in1;
  reg  [15:0] sram_out1;
  
  wire [15:0] sram_in2;
  reg  [15:0] sram_out2;
  
  wire [15:0] sram_in3;
  reg  [15:0] sram_out3;
  
  reg sram_wren0;
  reg sram_wren1;
  reg sram_wren2;
  reg sram_wren3;
 
  // SPRAM bank 0
 
      always @(posedge clk)
      begin
        if (io_wr & (mem_addr == `addr_sram_data0))
        begin
          sram_out0 <= dout;
          sram_wren0 <= 1;
        end else begin
          sram_wren0 <= 0;
        end
      end

    SB_SPRAM256KA  ramfn_inst0(
        .DATAIN(sram_out0),
        .ADDRESS(sram_addr),
        .MASKWREN(4'b1111),
        .WREN(sram_wren0),
        .CHIPSELECT(1'b1),
        .CLOCK(clk),
        .STANDBY(1'b0),
        .SLEEP(1'b0),
        .POWEROFF(1'b1),
        .DATAOUT(sram_in0)
);

  // SPRAM bank 1
 
      always @(posedge clk)
      begin
        if (io_wr & (mem_addr == `addr_sram_data1))
        begin
          sram_out1 <= dout;
          sram_wren1 <= 1;
        end else begin
          sram_wren1 <= 0;
        end
      end

    SB_SPRAM256KA  ramfn_inst1(
        .DATAIN(sram_out1),
        .ADDRESS(sram_addr),
        .MASKWREN(4'b1111),
        .WREN(sram_wren1),
        .CHIPSELECT(1'b1),
        .CLOCK(clk),
        .STANDBY(1'b0),
        .SLEEP(1'b0),
        .POWEROFF(1'b1),
        .DATAOUT(sram_in1)
    );

  // SPRAM bank 2
 
      always @(posedge clk)
      begin
        if (io_wr & (mem_addr == `addr_sram_data2))
        begin
          sram_out2 <= dout;
          sram_wren2 <= 1;
        end else begin
          sram_wren2 <= 0;
        end
      end

    SB_SPRAM256KA  ramfn_inst2(
        .DATAIN(sram_out2),
        .ADDRESS(sram_addr),
        .MASKWREN(4'b1111),
        .WREN(sram_wren2),
        .CHIPSELECT(1'b1),
        .CLOCK(clk),
        .STANDBY(1'b0),
        .SLEEP(1'b0),
        .POWEROFF(1'b1),
        .DATAOUT(sram_in2)
    );

  // SPRAM bank 3
 
      always @(posedge clk)
      begin
        if (io_wr & (mem_addr == `addr_sram_data3))
        begin
          sram_out3 <= dout;
          sram_wren3 <= 1;
        end else begin
          sram_wren3 <= 0;
        end
      end

    SB_SPRAM256KA  ramfn_inst3(
        .DATAIN(sram_out3),
        .ADDRESS(sram_addr),
        .MASKWREN(4'b1111),
        .WREN(sram_wren3),
        .CHIPSELECT(1'b1),
        .CLOCK(clk),
        .STANDBY(1'b0),
        .SLEEP(1'b0),
        .POWEROFF(1'b1),
        .DATAOUT(sram_in3)
    );

endmodule // top
